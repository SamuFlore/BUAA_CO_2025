`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:37:25 09/11/2025
// Design Name:   elevator
// Module Name:   E:/CO/ISE/ISE_Project/elevator/elevator_tb.v
// Project Name:  elevator
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: elevator
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module elevator_tb;

    // �����ź�
    reg [2:0] from;
    reg clk;
    reg reset;
    
    // ����ź�
    wire out;
    wire [2:0] cur_floor;
    wire direction;
    wire [2:0] request;
    
    // ʵ����������ģ��
    elevator uut (
        .from(from),
        .clk(clk),
        .reset(reset),
        .out(out),
        .cur_floor(cur_floor),
        .direction(direction),
        .request(request)
    );
    
    // ����10ns���ڵ�ʱ�ӣ���0ʱ�̿�ʼ������ת��
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 5ns��תһ�Σ�����10ns
    end
    
    // ���Լ���
    initial begin
        // ��ʼ״̬����������Ϊx��ȷ��ǰ5ns�ź�δ��ʼ��
        from = 3'bxxx;
        reset = 1'bx;
        
        // 5nsʱ����ʼ��ϵͳ�����ø�λ�ź�
        #5;
        reset = 1;         // ���λ
        from = 3'b000;     // ������
        
        // 15nsʱ���ͷŸ�λ��ȷ����λ����ά��һ��ʱ�����ڣ�
        #10;
        reset = 0;
        
        // 30nsʱ������1¥ָ���ǰʱ��=15+15=30ns��
        #15;
        from = 3'b001;     // 1¥����
        
        // 40nsʱ��ȡ������ά��һ��ʱ�����ڣ�
        #10;
        from = 3'b000;
        
        // 100nsʱ������5¥ָ���ǰʱ��=40+60=100ns��
        #60;
        from = 3'b101;     // 5¥����
        
        // 110nsʱ��ȡ������
        #10;
        from = 3'b000;
        
        // ��������һ��ʱ��۲���
        #200;
        
        // ��������

    end
    
endmodule
